module ModuloAnd(
   input IN0,
	input IN1,
	input IN2,
	input IN3,
	output OUT);
	
	assign OUT = IN0 & IN1 & IN2 & IN3;
	
endmodule
